`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 12/12/2018 02:03:19 AM
// Design Name: 
// Module Name: checkin
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module checkin(
    input [3:0] selector,
    input [10:0] timer,
    output reg [10:0] p1, p2, p3, p4 /* Parking check in time */
    );
   
    
endmodule
