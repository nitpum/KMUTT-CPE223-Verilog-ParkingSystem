`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 12/11/2018 05:30:53 PM
// Design Name: 
// Module Name: price_calculator
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module price_calculator(
    input enable,
    input [10:0] start_time, 
    input [10:0] end_time,
    input [6:0] price, // Max price 64
    output reg [17:0] value // Max value 1024 value = (end_time - start_time) / 60 * price
);
    always @ (posedge enable)
        begin
            if (enable)
                value <= (end_time - start_time) / 60 * price;
            else
                value = 0;
        end
endmodule
